module SQRT(

    input clk
    input [31:0] num;
    output sqrt;

    reg [31:0] a;
    reg [15:0] q;
    reg [17:0] left,right,r;

    integer i;
    
    );

    always_ff @(posedge clk)
        a = num;
        q = 0;
        i = 0;
        left = 0;   //input to adder/sub
        right = 0;  //input to adder/sub
        r = 0;  //remainder
        //run the calculations for 16 iterations.
        for(i=0;i<16;i=i+1) begin 
            right = {q,r[17],1'b1};
            left = {r[15:0],a[31:30]};
            a = {a[29:0],2'b00};    //left shift by 2 bits.
            if (r[17] == 1) //add if r is negative
                r = left + right;
            else    //subtract if r is positive
                r = left - right;
            q = {q[14:0],!r[17]};       
        end
        sqrt = q;   //final assignment of output.

    end

endmodule